`timescale 1ns / 1ps

module mousecontroler(
    );


endmodule
